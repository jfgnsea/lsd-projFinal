library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ROM_64_8 is
port(	address	:	in  std_logic_vector(5 downto 0);
		choiceBit:	in	 std_logic_vector;
		dataOut	:	out std_logic_vector(7 downto 0));
end ROM_64_8;

architecture Behavior of ROM_64_8 is

	type TROM is array (0 to 127) of std_logic_vector(7 downto 0); 
	-- valores aleatorios
	constant rom_mem: TROM := ("00101010", "11100111", "00010111", "10101000", "00010100", "01001110", "11010111", "11110000", 
										"00101011", "10110011", "10110100", "10111111", "01011011", "00001000", "01111001", "11110010", 
										"00001110", "00010010", "01001000", "00101000", "00011001", "00111001", "10011101", "01101011", 
										"10110101", "11000100", "10011001", "11011011", "11100101", "00001001", "10111010", "11111110", 
										"11010100", "10001001", "11111011", "01010001", "00010101", "01110101", "11111110", "00001010", 
										"00110011", "00010110", "11101101", "01000001", "00101101", "11001000", "10101000", "10010111", 
										"10110110", "11110100", "01110101", "01100011", "10101110", "00100001", "10100000", "10001110", 
										"10100010", "11010100", "11010101", "11000001", "10010011", "01001011", "01011101", "00111000",
										--segunda secçao da rom
										"11100001", "10011110", "01100010", "11011100", "00110101", "01111100", "00100001", "11011111", 
										"00000100", "11011110", "00000010", "01110100", "10100101", "10001011", "10001100", "01111010",
										"11100011", "01101010", "11100100", "00000001", "01000000", "00010100", "11010100", "01010111", 
										"00010100", "01110010", "00100100", "00000010", "00101001", "11011011", "01010111", "11011010", 
										"10110110", "11010001", "00101010", "10001111", "11000101", "00110010", "01001101", "01000111", 
										"00101110", "10000000", "01010111", "00111111", "11111110", "10111001", "11101001", "00011100", 
										"11001110", "11010000", "00101011", "01101100", "10000110", "10011010", "10111000", "11111110", 
										"11000001", "00000011", "10001110", "00001110", "00011111", "00101011", "01101010", "10111110"); 
	

begin

	dataOut <= rom_mem(to_integer(unsigned(choiceBit(0)&address)));

end Behavior;